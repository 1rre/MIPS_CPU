`timescale 1ps/1ps
module harvard_decode (
  
);

endmodule