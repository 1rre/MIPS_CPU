`timescale 1ps/1ps
module alu (
  input [31:0]
    a, b,
  output[31:0]
    r,
  output
    block
);



endmodule